top.sv
dut_interface.sv 
sequence_item.sv 
sequencer.sv 
sequence.sv 
subscriber.sv 
driver.sv  
monitor.sv
scoreboard.sv  
agent.sv
env.sv   
rsa_test.sv  
euclidean_loop.v  
gcd.v      
pt_exp.v     
RSA_decryptor.v        
encryption_key.v  
fifo.v            
lfsr.v     
multiply.v          
rsa_dut.sv         
RSA_encryptor.v                  
modexp1.v 
primality_tester.v  
 



 
